/*
	Emily Fredette
	request unit
*/

// interface
`include "request_unit_if.vh"

module request_unit (
  input CLK, nRST,
  request_unit_if.ru ruif
);

assign ruif.pcenable = ruif.ihit;

always_ff @(posedge CLK, negedge nRST) begin
	if (!nRST) begin
		ruif.dmemren = 0;
		ruif.dmemwen = 0;
	end
	else begin
		if (ruif.dhit) begin
			ruif.dmemren = 0;
			ruif.dmemwen = 0;
		end
		else begin
			//if (ruif.dwen) begin
			if (ruif.ihit & ruif.dwen) begin
				ruif.dmemwen = 1;
				ruif.dmemren = 0;
			end

			//if (ruif.dren) begin
			if (ruif.ihit & ruif.dren) begin
				ruif.dmemren = 1;
				ruif.dmemwen = 0;
			end
		end
	end
end

endmodule
