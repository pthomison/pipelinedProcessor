btb.sv
