/*
  Patrick Thomison
*/

// interface include
`include "cache_control_if.vh"

// memory types
`include "cpu_types_pkg.vh"

module dcache (
  input CLK, nRST,
  datapath_cache_if.cache dcif, 
  caches_if.caches cif
);

import cpu_types_pkg::*;

typedef struct packed {
	word_t wordA; 
	word_t wordB;
} block;

typedef struct packed {
	dcachef_t addr;
	block     data;
	logic     valid;
	logic     dirty
} frame;

frame cacheOne [15:0];
frame cacheTwo [15:0];

logic recUsed [15:0];

dcachef_t reqAddr, destCurrAddr;
word_t cdata, mload, mstore;

logic updateRead, updateWrite;

word_t loadAddrA, loadAddrB;

logic destination; // 0 for A, 1 for B

logic destinationDirty;

controllerState currState;
controllerState nextState;

typedef enum logic [3:0] {
IDLE         = 4'h0,
READHIT      = 4'h1,
MISSCHECK    = 4'h2,
WRITEHIT     = 4'h3,
DIRTYCLEANA  = 4'h4,
DIRTYCLEANB  = 4'h5,
READREQA     = 4'h6,
READREQB     = 4'h7,
READLOADA    = 4'h8,
READLOADB    = 4'h9,
FLUSH        = 4'hA,
STOP         = 4'hB
} controllerState;


// Type Casting To ICache Address
assign reqAddr = icachef_t'(dcif.imemaddr);

// Connecting mem data
assign mload   = cif.iload;
assign mstore  = dcif.dmemstore;

// Cache One Data Reg
// Handles nRST and writing in new values
always_ff @(posedge CLK, negedge nRST) begin
	if(nRST == 0) begin
		cacheOne    <= '{default:'0};
	end else begin
		if (destination == 0) begin
			if (updateRead == 1) begin
				cacheOne[reqAddr.idx].addr.tag    <= reqAddr.tag;
				cacheOne[reqAddr.idx].addr.idx    <= reqAddr.idx;
				cacheOne[reqAddr.idx].addr.bytoff <= reqAddr.bytoff;
				cacheOne[reqAddr.idx].data        <= mload;
				cacheOne[reqAddr.idx].valid       <= 1;
				cacheOne[reqAddr.idx].dirty       <= 0;
				recUsed[reqAddr.idx]              <= 0;
			end

			if (updateWrite == 1) begin
				cacheOne[reqAddr.idx].addr.tag    <= reqAddr.tag;
				cacheOne[reqAddr.idx].addr.idx    <= reqAddr.idx;
				cacheOne[reqAddr.idx].addr.bytoff <= reqAddr.bytoff;
				//cacheOne[reqAddr.idx].data        <= mstore;
				cacheOne[reqAddr.idx].valid       <= 1;
				cacheOne[reqAddr.idx].dirty       <= 1;

				if (reqAddr.blkoff == 0) begin
					cacheOne[reqAddr.idx].data.wordA <= mstore;
				end else begin
					cacheOne[reqAddr.idx].data.wordB <= mstore;
				end
			end
		end
	end
end

// Cache Two Data Reg
// Handles nRST and writing in new values
always_ff @(posedge CLK, negedge nRST) begin
	if(nRST == 0) begin
		cacheTwo    <= '{default:'0};
	end else begin
		if (destination == 1) begin
			if (updateRead == 1) begin
				cacheTwo[reqAddr.idx].addr.tag    <= reqAddr.tag;
				cacheTwo[reqAddr.idx].addr.idx    <= reqAddr.idx;
				cacheTwo[reqAddr.idx].addr.bytoff <= reqAddr.bytoff;
				cacheTwo[reqAddr.idx].data        <= mload;
				cacheTwo[reqAddr.idx].valid       <= 1;
				cacheTwo[reqAddr.idx].dirty       <= 0;
				recUsed[reqAddr.idx]              <= 1;
			end

			if (updateWrite == 1) begin
				cacheTwo[reqAddr.idx].addr.tag    <= reqAddr.tag;
				cacheTwo[reqAddr.idx].addr.idx    <= reqAddr.idx;
				cacheTwo[reqAddr.idx].addr.bytoff <= reqAddr.bytoff;
				cacheTwo[reqAddr.idx].data        <= mstore;
				cacheTwo[reqAddr.idx].valid       <= 1;
				cacheTwo[reqAddr.idx].dirty       <= 1;

				if (reqAddr.blkoff == 0) begin
					cacheTwo[reqAddr.idx].data.wordA <= mstore;
				end else begin
					cacheTwo[reqAddr.idx].data.wordB <= mstore;
				end
			end
		end
	end
end

// ----------------------------------------- //

assign prehitOne = (cacheOne[reqAddr.idx].addr.tag == reqAddr.tag) && (cacheOne[reqAddr.idx].valid == 1);
assign prehitTwo = (cacheTwo[reqAddr.idx].addr.tag == reqAddr.tag) && (cacheTwo[reqAddr.idx].valid == 1);
assign prehit = prehitOne || prehitTwo;

// ----------------------------------------- //

cdataOne = (reqAddr.blkoff == 0) ? cacheOne[reqAddr.idx].data.wordA : cacheOne[reqAddr.idx].data.wordB;
cdataTwo = (reqAddr.blkoff == 0) ? cacheTwo[reqAddr.idx].data.wordA : cacheTwo[reqAddr.idx].data.wordB;
cdata    = (prehitOne == 1) ? cdataOne : cdataTwo; // JANKY BAD TERRIBLE CODE; PLEASE FIX

// ----------------------------------------- //

// desination selector block
always_comb begin
	casez({validOne, validTwo})
		0: desination = 0;
		1: desination = 0;
		2: desination = 1;
		3: desination = (recentUsedOne == 1) 0 : 1;
		default: desination = 0;
	endcase

	if (desination == 0) begin
		dirtyAddr = cacheOne[reqAddr.idx].addr;
		dirtyData = cacheOne[reqAddr.idx].data;
	end else begin
		dirtyAddr = cacheTwo[reqAddr.idx].addr;
		dirtyData = cacheTwo[reqAddr.idx].data;
	end

	if (desination == 0) && (cacheOne[reqAddr.idx].dirty == 1) begin
		destinationDirty = 1;
	end else if (desination == 1) && (cacheTwo[reqAddr.idx].dirty == 1) begin
		destinationDirty = 1;
	end else begin
		destinationDirty = 0;
	end

end

// ----------------------------------------- //

// Determines correct address to request
always_comb begin
	if (reqAddr.blkoff == 0) begin
		loadAddrA = reqAddr.addr;
		loadAddrB = reqAddr.addr + 4;
	end else begin
		loadAddrA = reqAddr.addr - 4;
		loadAddrB = reqAddr.addr;
	end
end

// ----------------------------------------- //

// Cache Controller
// Handles nRST and advancing state
always_ff @(posedge CLK, negedge nRST) begin
	if(nRST == 0) begin
		currState <= IDLE;
	end else begin
		currState <= nextState;
	end
end

// Cache Controller
// Handles nextState and control signals
// Datapath Control Signals: dcif.dhit, dcif.dmemload, dcif.flushed
// RAM Control Signals: cif.dREN, cif.dWEN, cif.daddr, cif.dstore,
// Internal Control Signals: updateRead, updateWrite
always_comb begin
	if (currState == IDLE) begin
		dcif.dhit     = 0;
		dcif.dmemload = 0;
		dcif.flushed  = 0;

		cif.dREN      = 0;
		cif.dWEN      = 0;
		cif.daddr     = 0;
		cif.dstore    = 0;

		updateRead    = 0;
		updateWrite   = 0;

		if (dcif.halt == 1) begin
			nextState = FLUSH;

		end else if (dcif.dmemREN == 0 && dcif.dmemWEN == 0) begin
			nextState = IDLE;

		end else if (dcif.dmemREN == 1 && prehit == 1) begin
			// Read Hit;
			nextState = READHIT;

		end else if (dcif.dmemWEN == 1 && prehit == 1) begin
			// Write Hit;
			nextState = WRITEHIT;

		end else if (destinationDirty == 0) begin
			// Read Miss; Destination is NOT dirty
			nextState = READREQA;

		end else if (destinationDirty == 1) begin
			// Read Miss; Destination IS dirty
			nextState = DIRTYCLEANA;
		end

	end else if (currState == DIRTYCLEANA) begin
	// Writes Dirty Data (first word) Back To Memory

		dcif.dhit     = 0;
		dcif.dmemload = 0;
		dcif.flushed  = 0;

		cif.dREN      = 0;
		cif.dWEN      = 1;
		cif.daddr     = dirtyAddr;
		cif.dstore    = dirtyData.wordA;

		updateRead    = 0;
		updateWrite   = 0;

		if (cif.dwait == 1) begin
			nextState = DIRTYCLEANA;
		end else begin
			nextState = DIRTYCLEANB;
		end

	end else if (currState == DIRTYCLEANB) begin
	// Writes Dirty Data (second word) Back To Memory

		dcif.dhit     = 0;
		dcif.dmemload = 0;
		dcif.flushed  = 0;

		cif.dREN      = 0;
		cif.dWEN      = 1;
		cif.daddr     = dirtyAddr + 4;
		cif.dstore    = dirtyData.wordB;

		updateRead    = 0;
		updateWrite   = 0;

		if (cif.dwait == 1) begin
			nextState = DIRTYCLEANB;
		end else begin
			nextState = DATAREQA;
		end

	end else if (currState == DATAREQA) begin
	// Requests First Block of Data

		dcif.dhit     = 0;
		dcif.dmemload = 0;
		dcif.flushed  = 0;

		cif.dREN      = 1;
		cif.dWEN      = 0;
		cif.daddr     = loadAddrA;
		cif.dstore    = 0;

		updateRead    = 0;
		updateWrite   = 0;

		if (cif.dwait == 1) begin
			nextState = DATAREQA;
		end else begin
			nextState = DATALOADA;
		end

	end else if (currState == DATALOADA) begin
	// Loads First Block of Data into Cache

		dcif.dhit     = 0;
		dcif.dmemload = 0;
		dcif.flushed  = 0;

		cif.dREN      = 0;
		cif.dWEN      = 0;
		cif.daddr     = 0;
		cif.dstore    = 0;

		updateRead    = 1;
		updateWrite   = 0;

		nextState = DATAREQB;

	end else if (currState == DATAREQB) begin
	// Requests Second Block of Data

		dcif.dhit     = 0;
		dcif.dmemload = 0;
		dcif.flushed  = 0;

		cif.dREN      = 1;
		cif.dWEN      = 0;
		cif.daddr     = loadAddrB;
		cif.dstore    = 0;

		updateRead    = 0;
		updateWrite   = 0;

		if (cif.dwait == 1) begin
			nextState = DATAREQB;
		end else begin
			nextState = DATALOADB;
		end

	end else if (currState == DATALOADB) begin
	// Loads Second Block of Data into Cache

		dcif.dhit     = 0;
		dcif.dmemload = 0;
		dcif.flushed  = 0;

		cif.dREN      = 0;
		cif.dWEN      = 0;
		cif.daddr     = 0;
		cif.dstore    = 0;

		updateRead    = 1;

		updateWrite   = 0;

		nextState = IDLE;

	end else if (currState == READHIT) begin
	// Returns cached data to user

		dcif.dhit     = 1;
		dcif.dmemload = cdata;
		dcif.flushed  = 0;

		cif.dREN      = 0;
		cif.dWEN      = 0;
		cif.daddr     = 0;
		cif.dstore    = 0;

		updateRead    = 0;
		updateWrite   = 0;

		nextState = IDLE;

	end else if (currState == WRITEHIT) begin
	// Write user data to cache

		dcif.dhit     = 1;
		dcif.dmemload = 0;
		dcif.flushed  = 0;

		cif.dREN      = 0;
		cif.dWEN      = 0;
		cif.daddr     = 0;
		cif.dstore    = 0;

		updateRead    = 0;
		updateWrite   = 1;

		nextState = IDLE;


	end 
end