/*
Patrick Thomison
Emily Fredette
hazard unit
*/
`include "cpu_types_pkg.vh"


module hazard_unit (
  hazard_unit_if huif
);

  import cpu_types_pkg::*;

always_comb begin 




end //comb

endmodule